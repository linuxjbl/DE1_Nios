// nios2e.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2e (
		input  wire        clk_clk,                            //                         clk.clk
		output wire [27:0] decode0_external_connection_export, // decode0_external_connection.export
		output wire [27:0] decode1_external_connection_export, // decode1_external_connection.export
		output wire [27:0] decode2_external_connection_export, // decode2_external_connection.export
		output wire [27:0] decode3_external_connection_export, // decode3_external_connection.export
		output wire [27:0] decode4_external_connection_export, // decode4_external_connection.export
		output wire [27:0] decode5_external_connection_export, // decode5_external_connection.export
		output wire [27:0] decode6_external_connection_export, // decode6_external_connection.export
		output wire [27:0] decode7_external_connection_export, // decode7_external_connection.export
		output wire [7:0]  hex0_external_connection_export,    //    hex0_external_connection.export
		output wire [7:0]  hex1_external_connection_export,    //    hex1_external_connection.export
		output wire [7:0]  hex2_external_connection_export,    //    hex2_external_connection.export
		output wire [7:0]  hex3_external_connection_export,    //    hex3_external_connection.export
		output wire [7:0]  hex4_external_connection_export,    //    hex4_external_connection.export
		output wire [7:0]  hex5_external_connection_export,    //    hex5_external_connection.export
		output wire [27:0] period0_external_connection_export, // period0_external_connection.export
		output wire [27:0] period1_external_connection_export, // period1_external_connection.export
		output wire [27:0] period2_external_connection_export, // period2_external_connection.export
		output wire [27:0] period3_external_connection_export, // period3_external_connection.export
		output wire [27:0] period4_external_connection_export, // period4_external_connection.export
		output wire [27:0] period5_external_connection_export, // period5_external_connection.export
		output wire [27:0] period6_external_connection_export, // period6_external_connection.export
		output wire [27:0] period7_external_connection_export, // period7_external_connection.export
		input  wire [3:0]  push_external_connection_export,    //    push_external_connection.export
		input  wire        reset_reset_n                       //                       reset.reset_n
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [18:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_period0_s1_chipselect;                      // mm_interconnect_0:PERIOD0_s1_chipselect -> PERIOD0:chipselect
	wire  [31:0] mm_interconnect_0_period0_s1_readdata;                        // PERIOD0:readdata -> mm_interconnect_0:PERIOD0_s1_readdata
	wire   [1:0] mm_interconnect_0_period0_s1_address;                         // mm_interconnect_0:PERIOD0_s1_address -> PERIOD0:address
	wire         mm_interconnect_0_period0_s1_write;                           // mm_interconnect_0:PERIOD0_s1_write -> PERIOD0:write_n
	wire  [31:0] mm_interconnect_0_period0_s1_writedata;                       // mm_interconnect_0:PERIOD0_s1_writedata -> PERIOD0:writedata
	wire         mm_interconnect_0_decode0_s1_chipselect;                      // mm_interconnect_0:DECODE0_s1_chipselect -> DECODE0:chipselect
	wire  [31:0] mm_interconnect_0_decode0_s1_readdata;                        // DECODE0:readdata -> mm_interconnect_0:DECODE0_s1_readdata
	wire   [1:0] mm_interconnect_0_decode0_s1_address;                         // mm_interconnect_0:DECODE0_s1_address -> DECODE0:address
	wire         mm_interconnect_0_decode0_s1_write;                           // mm_interconnect_0:DECODE0_s1_write -> DECODE0:write_n
	wire  [31:0] mm_interconnect_0_decode0_s1_writedata;                       // mm_interconnect_0:DECODE0_s1_writedata -> DECODE0:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                         // mm_interconnect_0:HEX0_s1_chipselect -> HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                           // HEX0:readdata -> mm_interconnect_0:HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                            // mm_interconnect_0:HEX0_s1_address -> HEX0:address
	wire         mm_interconnect_0_hex0_s1_write;                              // mm_interconnect_0:HEX0_s1_write -> HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                          // mm_interconnect_0:HEX0_s1_writedata -> HEX0:writedata
	wire  [31:0] mm_interconnect_0_push_s1_readdata;                           // PUSH:readdata -> mm_interconnect_0:PUSH_s1_readdata
	wire   [1:0] mm_interconnect_0_push_s1_address;                            // mm_interconnect_0:PUSH_s1_address -> PUSH:address
	wire         mm_interconnect_0_period1_s1_chipselect;                      // mm_interconnect_0:PERIOD1_s1_chipselect -> PERIOD1:chipselect
	wire  [31:0] mm_interconnect_0_period1_s1_readdata;                        // PERIOD1:readdata -> mm_interconnect_0:PERIOD1_s1_readdata
	wire   [1:0] mm_interconnect_0_period1_s1_address;                         // mm_interconnect_0:PERIOD1_s1_address -> PERIOD1:address
	wire         mm_interconnect_0_period1_s1_write;                           // mm_interconnect_0:PERIOD1_s1_write -> PERIOD1:write_n
	wire  [31:0] mm_interconnect_0_period1_s1_writedata;                       // mm_interconnect_0:PERIOD1_s1_writedata -> PERIOD1:writedata
	wire         mm_interconnect_0_period2_s1_chipselect;                      // mm_interconnect_0:PERIOD2_s1_chipselect -> PERIOD2:chipselect
	wire  [31:0] mm_interconnect_0_period2_s1_readdata;                        // PERIOD2:readdata -> mm_interconnect_0:PERIOD2_s1_readdata
	wire   [1:0] mm_interconnect_0_period2_s1_address;                         // mm_interconnect_0:PERIOD2_s1_address -> PERIOD2:address
	wire         mm_interconnect_0_period2_s1_write;                           // mm_interconnect_0:PERIOD2_s1_write -> PERIOD2:write_n
	wire  [31:0] mm_interconnect_0_period2_s1_writedata;                       // mm_interconnect_0:PERIOD2_s1_writedata -> PERIOD2:writedata
	wire         mm_interconnect_0_period3_s1_chipselect;                      // mm_interconnect_0:PERIOD3_s1_chipselect -> PERIOD3:chipselect
	wire  [31:0] mm_interconnect_0_period3_s1_readdata;                        // PERIOD3:readdata -> mm_interconnect_0:PERIOD3_s1_readdata
	wire   [1:0] mm_interconnect_0_period3_s1_address;                         // mm_interconnect_0:PERIOD3_s1_address -> PERIOD3:address
	wire         mm_interconnect_0_period3_s1_write;                           // mm_interconnect_0:PERIOD3_s1_write -> PERIOD3:write_n
	wire  [31:0] mm_interconnect_0_period3_s1_writedata;                       // mm_interconnect_0:PERIOD3_s1_writedata -> PERIOD3:writedata
	wire         mm_interconnect_0_period4_s1_chipselect;                      // mm_interconnect_0:PERIOD4_s1_chipselect -> PERIOD4:chipselect
	wire  [31:0] mm_interconnect_0_period4_s1_readdata;                        // PERIOD4:readdata -> mm_interconnect_0:PERIOD4_s1_readdata
	wire   [1:0] mm_interconnect_0_period4_s1_address;                         // mm_interconnect_0:PERIOD4_s1_address -> PERIOD4:address
	wire         mm_interconnect_0_period4_s1_write;                           // mm_interconnect_0:PERIOD4_s1_write -> PERIOD4:write_n
	wire  [31:0] mm_interconnect_0_period4_s1_writedata;                       // mm_interconnect_0:PERIOD4_s1_writedata -> PERIOD4:writedata
	wire         mm_interconnect_0_period5_s1_chipselect;                      // mm_interconnect_0:PERIOD5_s1_chipselect -> PERIOD5:chipselect
	wire  [31:0] mm_interconnect_0_period5_s1_readdata;                        // PERIOD5:readdata -> mm_interconnect_0:PERIOD5_s1_readdata
	wire   [1:0] mm_interconnect_0_period5_s1_address;                         // mm_interconnect_0:PERIOD5_s1_address -> PERIOD5:address
	wire         mm_interconnect_0_period5_s1_write;                           // mm_interconnect_0:PERIOD5_s1_write -> PERIOD5:write_n
	wire  [31:0] mm_interconnect_0_period5_s1_writedata;                       // mm_interconnect_0:PERIOD5_s1_writedata -> PERIOD5:writedata
	wire         mm_interconnect_0_period6_s1_chipselect;                      // mm_interconnect_0:PERIOD6_s1_chipselect -> PERIOD6:chipselect
	wire  [31:0] mm_interconnect_0_period6_s1_readdata;                        // PERIOD6:readdata -> mm_interconnect_0:PERIOD6_s1_readdata
	wire   [1:0] mm_interconnect_0_period6_s1_address;                         // mm_interconnect_0:PERIOD6_s1_address -> PERIOD6:address
	wire         mm_interconnect_0_period6_s1_write;                           // mm_interconnect_0:PERIOD6_s1_write -> PERIOD6:write_n
	wire  [31:0] mm_interconnect_0_period6_s1_writedata;                       // mm_interconnect_0:PERIOD6_s1_writedata -> PERIOD6:writedata
	wire         mm_interconnect_0_period7_s1_chipselect;                      // mm_interconnect_0:PERIOD7_s1_chipselect -> PERIOD7:chipselect
	wire  [31:0] mm_interconnect_0_period7_s1_readdata;                        // PERIOD7:readdata -> mm_interconnect_0:PERIOD7_s1_readdata
	wire   [1:0] mm_interconnect_0_period7_s1_address;                         // mm_interconnect_0:PERIOD7_s1_address -> PERIOD7:address
	wire         mm_interconnect_0_period7_s1_write;                           // mm_interconnect_0:PERIOD7_s1_write -> PERIOD7:write_n
	wire  [31:0] mm_interconnect_0_period7_s1_writedata;                       // mm_interconnect_0:PERIOD7_s1_writedata -> PERIOD7:writedata
	wire         mm_interconnect_0_decode1_s1_chipselect;                      // mm_interconnect_0:DECODE1_s1_chipselect -> DECODE1:chipselect
	wire  [31:0] mm_interconnect_0_decode1_s1_readdata;                        // DECODE1:readdata -> mm_interconnect_0:DECODE1_s1_readdata
	wire   [1:0] mm_interconnect_0_decode1_s1_address;                         // mm_interconnect_0:DECODE1_s1_address -> DECODE1:address
	wire         mm_interconnect_0_decode1_s1_write;                           // mm_interconnect_0:DECODE1_s1_write -> DECODE1:write_n
	wire  [31:0] mm_interconnect_0_decode1_s1_writedata;                       // mm_interconnect_0:DECODE1_s1_writedata -> DECODE1:writedata
	wire         mm_interconnect_0_decode2_s1_chipselect;                      // mm_interconnect_0:DECODE2_s1_chipselect -> DECODE2:chipselect
	wire  [31:0] mm_interconnect_0_decode2_s1_readdata;                        // DECODE2:readdata -> mm_interconnect_0:DECODE2_s1_readdata
	wire   [1:0] mm_interconnect_0_decode2_s1_address;                         // mm_interconnect_0:DECODE2_s1_address -> DECODE2:address
	wire         mm_interconnect_0_decode2_s1_write;                           // mm_interconnect_0:DECODE2_s1_write -> DECODE2:write_n
	wire  [31:0] mm_interconnect_0_decode2_s1_writedata;                       // mm_interconnect_0:DECODE2_s1_writedata -> DECODE2:writedata
	wire         mm_interconnect_0_decode3_s1_chipselect;                      // mm_interconnect_0:DECODE3_s1_chipselect -> DECODE3:chipselect
	wire  [31:0] mm_interconnect_0_decode3_s1_readdata;                        // DECODE3:readdata -> mm_interconnect_0:DECODE3_s1_readdata
	wire   [1:0] mm_interconnect_0_decode3_s1_address;                         // mm_interconnect_0:DECODE3_s1_address -> DECODE3:address
	wire         mm_interconnect_0_decode3_s1_write;                           // mm_interconnect_0:DECODE3_s1_write -> DECODE3:write_n
	wire  [31:0] mm_interconnect_0_decode3_s1_writedata;                       // mm_interconnect_0:DECODE3_s1_writedata -> DECODE3:writedata
	wire         mm_interconnect_0_decode4_s1_chipselect;                      // mm_interconnect_0:DECODE4_s1_chipselect -> DECODE4:chipselect
	wire  [31:0] mm_interconnect_0_decode4_s1_readdata;                        // DECODE4:readdata -> mm_interconnect_0:DECODE4_s1_readdata
	wire   [1:0] mm_interconnect_0_decode4_s1_address;                         // mm_interconnect_0:DECODE4_s1_address -> DECODE4:address
	wire         mm_interconnect_0_decode4_s1_write;                           // mm_interconnect_0:DECODE4_s1_write -> DECODE4:write_n
	wire  [31:0] mm_interconnect_0_decode4_s1_writedata;                       // mm_interconnect_0:DECODE4_s1_writedata -> DECODE4:writedata
	wire         mm_interconnect_0_decode5_s1_chipselect;                      // mm_interconnect_0:DECODE5_s1_chipselect -> DECODE5:chipselect
	wire  [31:0] mm_interconnect_0_decode5_s1_readdata;                        // DECODE5:readdata -> mm_interconnect_0:DECODE5_s1_readdata
	wire   [1:0] mm_interconnect_0_decode5_s1_address;                         // mm_interconnect_0:DECODE5_s1_address -> DECODE5:address
	wire         mm_interconnect_0_decode5_s1_write;                           // mm_interconnect_0:DECODE5_s1_write -> DECODE5:write_n
	wire  [31:0] mm_interconnect_0_decode5_s1_writedata;                       // mm_interconnect_0:DECODE5_s1_writedata -> DECODE5:writedata
	wire         mm_interconnect_0_decode6_s1_chipselect;                      // mm_interconnect_0:DECODE6_s1_chipselect -> DECODE6:chipselect
	wire  [31:0] mm_interconnect_0_decode6_s1_readdata;                        // DECODE6:readdata -> mm_interconnect_0:DECODE6_s1_readdata
	wire   [1:0] mm_interconnect_0_decode6_s1_address;                         // mm_interconnect_0:DECODE6_s1_address -> DECODE6:address
	wire         mm_interconnect_0_decode6_s1_write;                           // mm_interconnect_0:DECODE6_s1_write -> DECODE6:write_n
	wire  [31:0] mm_interconnect_0_decode6_s1_writedata;                       // mm_interconnect_0:DECODE6_s1_writedata -> DECODE6:writedata
	wire         mm_interconnect_0_decode7_s1_chipselect;                      // mm_interconnect_0:DECODE7_s1_chipselect -> DECODE7:chipselect
	wire  [31:0] mm_interconnect_0_decode7_s1_readdata;                        // DECODE7:readdata -> mm_interconnect_0:DECODE7_s1_readdata
	wire   [1:0] mm_interconnect_0_decode7_s1_address;                         // mm_interconnect_0:DECODE7_s1_address -> DECODE7:address
	wire         mm_interconnect_0_decode7_s1_write;                           // mm_interconnect_0:DECODE7_s1_write -> DECODE7:write_n
	wire  [31:0] mm_interconnect_0_decode7_s1_writedata;                       // mm_interconnect_0:DECODE7_s1_writedata -> DECODE7:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                         // mm_interconnect_0:HEX1_s1_chipselect -> HEX1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                           // HEX1:readdata -> mm_interconnect_0:HEX1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                            // mm_interconnect_0:HEX1_s1_address -> HEX1:address
	wire         mm_interconnect_0_hex1_s1_write;                              // mm_interconnect_0:HEX1_s1_write -> HEX1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                          // mm_interconnect_0:HEX1_s1_writedata -> HEX1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                         // mm_interconnect_0:HEX2_s1_chipselect -> HEX2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                           // HEX2:readdata -> mm_interconnect_0:HEX2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                            // mm_interconnect_0:HEX2_s1_address -> HEX2:address
	wire         mm_interconnect_0_hex2_s1_write;                              // mm_interconnect_0:HEX2_s1_write -> HEX2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                          // mm_interconnect_0:HEX2_s1_writedata -> HEX2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                         // mm_interconnect_0:HEX3_s1_chipselect -> HEX3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                           // HEX3:readdata -> mm_interconnect_0:HEX3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                            // mm_interconnect_0:HEX3_s1_address -> HEX3:address
	wire         mm_interconnect_0_hex3_s1_write;                              // mm_interconnect_0:HEX3_s1_write -> HEX3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                          // mm_interconnect_0:HEX3_s1_writedata -> HEX3:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                         // mm_interconnect_0:HEX4_s1_chipselect -> HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                           // HEX4:readdata -> mm_interconnect_0:HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                            // mm_interconnect_0:HEX4_s1_address -> HEX4:address
	wire         mm_interconnect_0_hex4_s1_write;                              // mm_interconnect_0:HEX4_s1_write -> HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                          // mm_interconnect_0:HEX4_s1_writedata -> HEX4:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                         // mm_interconnect_0:HEX5_s1_chipselect -> HEX5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                           // HEX5:readdata -> mm_interconnect_0:HEX5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                            // mm_interconnect_0:HEX5_s1_address -> HEX5:address
	wire         mm_interconnect_0_hex5_s1_write;                              // mm_interconnect_0:HEX5_s1_write -> HEX5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                          // mm_interconnect_0:HEX5_s1_writedata -> HEX5:writedata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [DECODE0:reset_n, DECODE1:reset_n, DECODE2:reset_n, DECODE3:reset_n, DECODE4:reset_n, DECODE5:reset_n, DECODE6:reset_n, DECODE7:reset_n, HEX0:reset_n, HEX1:reset_n, HEX2:reset_n, HEX3:reset_n, HEX4:reset_n, HEX5:reset_n, PERIOD0:reset_n, PERIOD1:reset_n, PERIOD2:reset_n, PERIOD3:reset_n, PERIOD4:reset_n, PERIOD5:reset_n, PERIOD6:reset_n, PERIOD7:reset_n, PUSH:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios2e_DECODE0 decode0 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode0_s1_readdata),   //                    .readdata
		.out_port   (decode0_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode1_s1_readdata),   //                    .readdata
		.out_port   (decode1_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode2_s1_readdata),   //                    .readdata
		.out_port   (decode2_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode3_s1_readdata),   //                    .readdata
		.out_port   (decode3_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode4 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode4_s1_readdata),   //                    .readdata
		.out_port   (decode4_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode5 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode5_s1_readdata),   //                    .readdata
		.out_port   (decode5_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode6 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode6_s1_readdata),   //                    .readdata
		.out_port   (decode6_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 decode7 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_decode7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_decode7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_decode7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_decode7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_decode7_s1_readdata),   //                    .readdata
		.out_port   (decode7_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_external_connection_export)       // external_connection.export
	);

	nios2e_HEX0 hex5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period0 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period0_s1_readdata),   //                    .readdata
		.out_port   (period0_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period1_s1_readdata),   //                    .readdata
		.out_port   (period1_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period2_s1_readdata),   //                    .readdata
		.out_port   (period2_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period3_s1_readdata),   //                    .readdata
		.out_port   (period3_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period4 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period4_s1_readdata),   //                    .readdata
		.out_port   (period4_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period5 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period5_s1_readdata),   //                    .readdata
		.out_port   (period5_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period6 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period6_s1_readdata),   //                    .readdata
		.out_port   (period6_external_connection_export)       // external_connection.export
	);

	nios2e_DECODE0 period7 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_period7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_period7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_period7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_period7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_period7_s1_readdata),   //                    .readdata
		.out_port   (period7_external_connection_export)       // external_connection.export
	);

	nios2e_PUSH push (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_push_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_push_s1_readdata), //                    .readdata
		.in_port  (push_external_connection_export)     // external_connection.export
	);

	nios2e_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios2e_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios2e_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios2e_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.DECODE0_s1_address                               (mm_interconnect_0_decode0_s1_address),                         //                                 DECODE0_s1.address
		.DECODE0_s1_write                                 (mm_interconnect_0_decode0_s1_write),                           //                                           .write
		.DECODE0_s1_readdata                              (mm_interconnect_0_decode0_s1_readdata),                        //                                           .readdata
		.DECODE0_s1_writedata                             (mm_interconnect_0_decode0_s1_writedata),                       //                                           .writedata
		.DECODE0_s1_chipselect                            (mm_interconnect_0_decode0_s1_chipselect),                      //                                           .chipselect
		.DECODE1_s1_address                               (mm_interconnect_0_decode1_s1_address),                         //                                 DECODE1_s1.address
		.DECODE1_s1_write                                 (mm_interconnect_0_decode1_s1_write),                           //                                           .write
		.DECODE1_s1_readdata                              (mm_interconnect_0_decode1_s1_readdata),                        //                                           .readdata
		.DECODE1_s1_writedata                             (mm_interconnect_0_decode1_s1_writedata),                       //                                           .writedata
		.DECODE1_s1_chipselect                            (mm_interconnect_0_decode1_s1_chipselect),                      //                                           .chipselect
		.DECODE2_s1_address                               (mm_interconnect_0_decode2_s1_address),                         //                                 DECODE2_s1.address
		.DECODE2_s1_write                                 (mm_interconnect_0_decode2_s1_write),                           //                                           .write
		.DECODE2_s1_readdata                              (mm_interconnect_0_decode2_s1_readdata),                        //                                           .readdata
		.DECODE2_s1_writedata                             (mm_interconnect_0_decode2_s1_writedata),                       //                                           .writedata
		.DECODE2_s1_chipselect                            (mm_interconnect_0_decode2_s1_chipselect),                      //                                           .chipselect
		.DECODE3_s1_address                               (mm_interconnect_0_decode3_s1_address),                         //                                 DECODE3_s1.address
		.DECODE3_s1_write                                 (mm_interconnect_0_decode3_s1_write),                           //                                           .write
		.DECODE3_s1_readdata                              (mm_interconnect_0_decode3_s1_readdata),                        //                                           .readdata
		.DECODE3_s1_writedata                             (mm_interconnect_0_decode3_s1_writedata),                       //                                           .writedata
		.DECODE3_s1_chipselect                            (mm_interconnect_0_decode3_s1_chipselect),                      //                                           .chipselect
		.DECODE4_s1_address                               (mm_interconnect_0_decode4_s1_address),                         //                                 DECODE4_s1.address
		.DECODE4_s1_write                                 (mm_interconnect_0_decode4_s1_write),                           //                                           .write
		.DECODE4_s1_readdata                              (mm_interconnect_0_decode4_s1_readdata),                        //                                           .readdata
		.DECODE4_s1_writedata                             (mm_interconnect_0_decode4_s1_writedata),                       //                                           .writedata
		.DECODE4_s1_chipselect                            (mm_interconnect_0_decode4_s1_chipselect),                      //                                           .chipselect
		.DECODE5_s1_address                               (mm_interconnect_0_decode5_s1_address),                         //                                 DECODE5_s1.address
		.DECODE5_s1_write                                 (mm_interconnect_0_decode5_s1_write),                           //                                           .write
		.DECODE5_s1_readdata                              (mm_interconnect_0_decode5_s1_readdata),                        //                                           .readdata
		.DECODE5_s1_writedata                             (mm_interconnect_0_decode5_s1_writedata),                       //                                           .writedata
		.DECODE5_s1_chipselect                            (mm_interconnect_0_decode5_s1_chipselect),                      //                                           .chipselect
		.DECODE6_s1_address                               (mm_interconnect_0_decode6_s1_address),                         //                                 DECODE6_s1.address
		.DECODE6_s1_write                                 (mm_interconnect_0_decode6_s1_write),                           //                                           .write
		.DECODE6_s1_readdata                              (mm_interconnect_0_decode6_s1_readdata),                        //                                           .readdata
		.DECODE6_s1_writedata                             (mm_interconnect_0_decode6_s1_writedata),                       //                                           .writedata
		.DECODE6_s1_chipselect                            (mm_interconnect_0_decode6_s1_chipselect),                      //                                           .chipselect
		.DECODE7_s1_address                               (mm_interconnect_0_decode7_s1_address),                         //                                 DECODE7_s1.address
		.DECODE7_s1_write                                 (mm_interconnect_0_decode7_s1_write),                           //                                           .write
		.DECODE7_s1_readdata                              (mm_interconnect_0_decode7_s1_readdata),                        //                                           .readdata
		.DECODE7_s1_writedata                             (mm_interconnect_0_decode7_s1_writedata),                       //                                           .writedata
		.DECODE7_s1_chipselect                            (mm_interconnect_0_decode7_s1_chipselect),                      //                                           .chipselect
		.HEX0_s1_address                                  (mm_interconnect_0_hex0_s1_address),                            //                                    HEX0_s1.address
		.HEX0_s1_write                                    (mm_interconnect_0_hex0_s1_write),                              //                                           .write
		.HEX0_s1_readdata                                 (mm_interconnect_0_hex0_s1_readdata),                           //                                           .readdata
		.HEX0_s1_writedata                                (mm_interconnect_0_hex0_s1_writedata),                          //                                           .writedata
		.HEX0_s1_chipselect                               (mm_interconnect_0_hex0_s1_chipselect),                         //                                           .chipselect
		.HEX1_s1_address                                  (mm_interconnect_0_hex1_s1_address),                            //                                    HEX1_s1.address
		.HEX1_s1_write                                    (mm_interconnect_0_hex1_s1_write),                              //                                           .write
		.HEX1_s1_readdata                                 (mm_interconnect_0_hex1_s1_readdata),                           //                                           .readdata
		.HEX1_s1_writedata                                (mm_interconnect_0_hex1_s1_writedata),                          //                                           .writedata
		.HEX1_s1_chipselect                               (mm_interconnect_0_hex1_s1_chipselect),                         //                                           .chipselect
		.HEX2_s1_address                                  (mm_interconnect_0_hex2_s1_address),                            //                                    HEX2_s1.address
		.HEX2_s1_write                                    (mm_interconnect_0_hex2_s1_write),                              //                                           .write
		.HEX2_s1_readdata                                 (mm_interconnect_0_hex2_s1_readdata),                           //                                           .readdata
		.HEX2_s1_writedata                                (mm_interconnect_0_hex2_s1_writedata),                          //                                           .writedata
		.HEX2_s1_chipselect                               (mm_interconnect_0_hex2_s1_chipselect),                         //                                           .chipselect
		.HEX3_s1_address                                  (mm_interconnect_0_hex3_s1_address),                            //                                    HEX3_s1.address
		.HEX3_s1_write                                    (mm_interconnect_0_hex3_s1_write),                              //                                           .write
		.HEX3_s1_readdata                                 (mm_interconnect_0_hex3_s1_readdata),                           //                                           .readdata
		.HEX3_s1_writedata                                (mm_interconnect_0_hex3_s1_writedata),                          //                                           .writedata
		.HEX3_s1_chipselect                               (mm_interconnect_0_hex3_s1_chipselect),                         //                                           .chipselect
		.HEX4_s1_address                                  (mm_interconnect_0_hex4_s1_address),                            //                                    HEX4_s1.address
		.HEX4_s1_write                                    (mm_interconnect_0_hex4_s1_write),                              //                                           .write
		.HEX4_s1_readdata                                 (mm_interconnect_0_hex4_s1_readdata),                           //                                           .readdata
		.HEX4_s1_writedata                                (mm_interconnect_0_hex4_s1_writedata),                          //                                           .writedata
		.HEX4_s1_chipselect                               (mm_interconnect_0_hex4_s1_chipselect),                         //                                           .chipselect
		.HEX5_s1_address                                  (mm_interconnect_0_hex5_s1_address),                            //                                    HEX5_s1.address
		.HEX5_s1_write                                    (mm_interconnect_0_hex5_s1_write),                              //                                           .write
		.HEX5_s1_readdata                                 (mm_interconnect_0_hex5_s1_readdata),                           //                                           .readdata
		.HEX5_s1_writedata                                (mm_interconnect_0_hex5_s1_writedata),                          //                                           .writedata
		.HEX5_s1_chipselect                               (mm_interconnect_0_hex5_s1_chipselect),                         //                                           .chipselect
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.PERIOD0_s1_address                               (mm_interconnect_0_period0_s1_address),                         //                                 PERIOD0_s1.address
		.PERIOD0_s1_write                                 (mm_interconnect_0_period0_s1_write),                           //                                           .write
		.PERIOD0_s1_readdata                              (mm_interconnect_0_period0_s1_readdata),                        //                                           .readdata
		.PERIOD0_s1_writedata                             (mm_interconnect_0_period0_s1_writedata),                       //                                           .writedata
		.PERIOD0_s1_chipselect                            (mm_interconnect_0_period0_s1_chipselect),                      //                                           .chipselect
		.PERIOD1_s1_address                               (mm_interconnect_0_period1_s1_address),                         //                                 PERIOD1_s1.address
		.PERIOD1_s1_write                                 (mm_interconnect_0_period1_s1_write),                           //                                           .write
		.PERIOD1_s1_readdata                              (mm_interconnect_0_period1_s1_readdata),                        //                                           .readdata
		.PERIOD1_s1_writedata                             (mm_interconnect_0_period1_s1_writedata),                       //                                           .writedata
		.PERIOD1_s1_chipselect                            (mm_interconnect_0_period1_s1_chipselect),                      //                                           .chipselect
		.PERIOD2_s1_address                               (mm_interconnect_0_period2_s1_address),                         //                                 PERIOD2_s1.address
		.PERIOD2_s1_write                                 (mm_interconnect_0_period2_s1_write),                           //                                           .write
		.PERIOD2_s1_readdata                              (mm_interconnect_0_period2_s1_readdata),                        //                                           .readdata
		.PERIOD2_s1_writedata                             (mm_interconnect_0_period2_s1_writedata),                       //                                           .writedata
		.PERIOD2_s1_chipselect                            (mm_interconnect_0_period2_s1_chipselect),                      //                                           .chipselect
		.PERIOD3_s1_address                               (mm_interconnect_0_period3_s1_address),                         //                                 PERIOD3_s1.address
		.PERIOD3_s1_write                                 (mm_interconnect_0_period3_s1_write),                           //                                           .write
		.PERIOD3_s1_readdata                              (mm_interconnect_0_period3_s1_readdata),                        //                                           .readdata
		.PERIOD3_s1_writedata                             (mm_interconnect_0_period3_s1_writedata),                       //                                           .writedata
		.PERIOD3_s1_chipselect                            (mm_interconnect_0_period3_s1_chipselect),                      //                                           .chipselect
		.PERIOD4_s1_address                               (mm_interconnect_0_period4_s1_address),                         //                                 PERIOD4_s1.address
		.PERIOD4_s1_write                                 (mm_interconnect_0_period4_s1_write),                           //                                           .write
		.PERIOD4_s1_readdata                              (mm_interconnect_0_period4_s1_readdata),                        //                                           .readdata
		.PERIOD4_s1_writedata                             (mm_interconnect_0_period4_s1_writedata),                       //                                           .writedata
		.PERIOD4_s1_chipselect                            (mm_interconnect_0_period4_s1_chipselect),                      //                                           .chipselect
		.PERIOD5_s1_address                               (mm_interconnect_0_period5_s1_address),                         //                                 PERIOD5_s1.address
		.PERIOD5_s1_write                                 (mm_interconnect_0_period5_s1_write),                           //                                           .write
		.PERIOD5_s1_readdata                              (mm_interconnect_0_period5_s1_readdata),                        //                                           .readdata
		.PERIOD5_s1_writedata                             (mm_interconnect_0_period5_s1_writedata),                       //                                           .writedata
		.PERIOD5_s1_chipselect                            (mm_interconnect_0_period5_s1_chipselect),                      //                                           .chipselect
		.PERIOD6_s1_address                               (mm_interconnect_0_period6_s1_address),                         //                                 PERIOD6_s1.address
		.PERIOD6_s1_write                                 (mm_interconnect_0_period6_s1_write),                           //                                           .write
		.PERIOD6_s1_readdata                              (mm_interconnect_0_period6_s1_readdata),                        //                                           .readdata
		.PERIOD6_s1_writedata                             (mm_interconnect_0_period6_s1_writedata),                       //                                           .writedata
		.PERIOD6_s1_chipselect                            (mm_interconnect_0_period6_s1_chipselect),                      //                                           .chipselect
		.PERIOD7_s1_address                               (mm_interconnect_0_period7_s1_address),                         //                                 PERIOD7_s1.address
		.PERIOD7_s1_write                                 (mm_interconnect_0_period7_s1_write),                           //                                           .write
		.PERIOD7_s1_readdata                              (mm_interconnect_0_period7_s1_readdata),                        //                                           .readdata
		.PERIOD7_s1_writedata                             (mm_interconnect_0_period7_s1_writedata),                       //                                           .writedata
		.PERIOD7_s1_chipselect                            (mm_interconnect_0_period7_s1_chipselect),                      //                                           .chipselect
		.PUSH_s1_address                                  (mm_interconnect_0_push_s1_address),                            //                                    PUSH_s1.address
		.PUSH_s1_readdata                                 (mm_interconnect_0_push_s1_readdata)                            //                                           .readdata
	);

	nios2e_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
